module led(
  output blue_led
);

  assign blue_led = 0;

endmodule

