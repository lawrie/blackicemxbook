module rgbled(
	input [2:0] switch,
	output [2:0] rgb
);
	
	assign rgb = switch;
	
endmodule

