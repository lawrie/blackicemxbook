module led(
  output reg blue_led
);

  always @(*) blue_led = 0;

endmodule

