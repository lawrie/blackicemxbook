module button_test(
  output yellow_led,
  input button1
);

  assign yellow_led = button1;

endmodule

