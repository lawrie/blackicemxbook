module leds(
  output [3:0] leds
);

  assign leds = 4'b0000;

endmodule

